190020039 Dhruv Shah bjt_current_mirror

.SUBCKT ZENER_12 1 2 
D1 1 2 DF 
DZ 3 1 DR 
VZ 2 3 10.8 
.MODEL DF D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330 TT=50.1n ) 
.MODEL DR D ( IS=5.49f RS=50 N=1.77 ) 
.ENDS 
v1 1 0 12 
r1 1 2 10k 
Q1 2 2 0 bc547a 
Q2 4 2 0 bc547a 
v2 4 0 dc 1 ac 0 
.dc v2 1 5 0.5 

.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3  
+ BR=9.5 VAF=100 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40  
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f 

.control 
run 
print i(v2) 
.endc 
.end
