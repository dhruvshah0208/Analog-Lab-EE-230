skip-line

.SUBCKT ZENER_12 1 2
D1 1 2 DF
DZ 3 1 DR
VZ 2 3 10.8
.MODEL DF D ( IS=27.5p RS=0.620 N=1.10 CJO=78.3p VJ=1.00 M=0.330 TT=50.1n )
.MODEL DR D ( IS=5.49f RS=125 N=1.77 )
.ENDS

Vin in 0 20
Rs in dummy_r 470
vrdummy dummy_r out dc 0

vzdummy out dummy_z dc 0
x_zener 0 dummy_z ZENER_12

Rl out dummy_load 0
voutdummy dummy_load 0 dc 0

.dc Rl 100 1000 5
.control

run

plot v(in) v(out)
plot i(voutdummy) i(vrdummy) i(vzdummy)

.endc
.end
