Dhruv Shah 190020039
.model 1N4007 D (IS=5.44e-7 N=2.337 RS=0.0429 BV=1000 IBV=5u tnom=25e0)

v A B sin(0 21.213 50 1n 1n 1n)

D1 A dummy1 1N4007
vdummy1 dummy1 out dc 0

D2 B dummy3 1N4007
vdummy3 dummy3 out dc 0

D3 gnd A 1N4007

D4 gnd B 1N4007
Rl out gnd 1000
C out gnd 1000u

.tran 0.001 0.1

.control

run

plot i(vdummy1) i(vdummy3)
plot v(out)

set hcopydevtype=postscript
set hcopypscolor=1
hardcopy q1_plot1.ps i(vdummy1) i(vdummy3)
hardcopy q1_-plot2.ps v(out)

.endc
.end
