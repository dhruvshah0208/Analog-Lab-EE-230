Unregulated DC Power supply

.model 1N4007 D (IS=5.44e-7 N=2.337 RS=0.0429 BV=1000 IBV=5u tnom=25e0)
 
*.MODEL 1N914 D (IS=6.2229E-9  N=1.9224  RS=0.33636  IKF=42.843E-3  CJO=764.38E-15 
+ M=0.1001 VJ=0.99900  BV=100.14  IBV=0.25951  TT=2.8854E-9)

v A B sin(0 21.213 50)

D1 A dummy1 1N4007
vdummy1 dummy1 out dc 0

D2 B out 1N4007

D3 gnd dummy2 1N4007
vdummy2 dummy2 A dc 0

D4 gnd B 1N4007
Rl out gnd 1000

.tran 0.001 0.1

.control

run

set hcopydevtype=postscript
set hcopypscolor=1
*hardcopy unreg_currents.eps i(vdummy1) i(vdummy2)

plot i(vdummy1) i(vdummy2) v(out)
*plot v(A)-v(B)-v(out)

.endc
.end
