Dhruv Shah 190020039 RC Differentiator Circuit
*Circuit Description
r1 2 0 10k
c1 1 2 0.1u
*Voltage Description 
*v1n 1 0 pulse(0 5 delay rise_time fall_time T Period)
v1n 1 0 pulse(0 5 0 0 0 0.1m 0.2m)

*transient Analysis
*.tran step 3*periodz

.tran 0.01m 4m
.control
run

*Plotting
plot v(1) v(2)
set hcopypscolor = 1
hardcopy diff_final_pt1.ps v(1) v(2)
.endc
.end
