190020039 Dhruv Shah bjt_diff_amp

vcc 1 0 12 
rc1 1 17 6.8k 
rc2 1 18 6.8k 
vc1 17 2 0 
vc2 18 3 0 
Q1 2 5 4 bc547a 
Q2 3 6 4 bc547a 
re 4 7 10k 
vee 7 0 -12 
rb1 5 12 1k 
rb2 6 13 1k 
vin1 12 0 sin(0 10m 1k 0 0) 
vin2 13 0 0 
.tran
.model bc547a NPN IS=10f BF=200 ISE=10.3f IKF=50m NE=1.3  
+ BR=9.5 VAF=80 IKR=12m ISC=47p NC=2 VAR=10 RB=280 RE=1 RC=40  
+ tr=0.3u tf=0.5n cje=12p vje=0.48 mje=0.5 cjc=6p vjc=0.7 mjc=0.33 kf=2f 

.control 
run 
plot v(2) v(3)

.endc 
.end 
